package tb_global_mem_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh";
  `include "../tb_common/mat_conv.svh";
  `include "tb_global_mem_lsram_wrapper.svh";
  `include "tb_global_mem_usram_wrapper.svh";

endpackage
