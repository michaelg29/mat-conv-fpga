
`include "uvm_macros.svh"

import uvm_pkg::*;

// testcase exercising valid kernel command and payload
class tb_cluster_kernel_size_subject_no_pad 
  #(int KERNEL_SIZE = 5, 
    int FIFO_WIDTH = 8,
    int NUM_ROWS = 5,
    int NUM_COLS = 5) 
    extends mat_conv_tc;

  // virtual interfacepixel
  virtual cluster_if vif;

  // clock period definition
  time MACCLK_PER;

  int num_additional_cycles_shifts;

   // local params
  localparam PADDING = (KERNEL_SIZE-1)/2;

  // constructor
  function new(virtual cluster_if vif, time MACCLK_PER);
    this.vif = vif;
    this.MACCLK_PER = MACCLK_PER;
  endfunction // new

  task automatic run;
    //UNRESOLVED
    //logic [vif.KERNEL_SIZE-1:0][vif.KERNEL_SIZE-1:0][7:0] kernel;
    //logic [vif.KERNEL_SIZE-1:0][vif.KERNEL_SIZE-1:0][7:0] image;
    logic [KERNEL_SIZE-1:0][KERNEL_SIZE-1:0][7:0] kernel;
    logic [NUM_ROWS-1:0][NUM_COLS-1:0][7:0] image;
    logic [NUM_ROWS-2*PADDING-1:0][NUM_COLS-2*PADDING-1:0][7:0] imconv;

    logic sign = 1'b0;

    `uvm_info("tb_cluster_kernel_size_subject_no_pad", "Executing testcase", UVM_NONE);

    @(posedge vif.i_clk);

    // Generate kernel and load it
    kernel = vif.kernel_gen();
    vif.load_kernel(kernel, sign);

    // Generate image
    image = vif.image_gen_nopad();

    //Calculate convolution result (unsigned)
    imconv = vif.image_conv_nopad(image, kernel, sign);

    vif.display_conv_nopad(image, kernel, imconv);


    @(posedge vif.i_clk);

    vif.i_discont <= 1;
    vif.i_waddr <= 0;

    //Change values on falling edge (problems when doing rising edge)
    @(negedge vif.i_clk);

    vif.i_is_subj <= 1;
    for (int row = 0 ; row < NUM_ROWS ; row++) begin
      vif.i_newrow <= 1;
      for (int col = 0 ; col < NUM_COLS ; col+=FIFO_WIDTH) begin
        vif.i_new_pkt <= 1;
        vif.i_pkt <= image[row][col +: FIFO_WIDTH]; //args must be multiple of FIFO_WIDTH
        
        @(negedge vif.i_clk);
        vif.i_newrow <= 0;

        //Image size is assumed to be a multiple of 128 (FIFO_WIDTH aligned). Always an additional 3 clock cycles delay
        num_additional_cycles_shifts = FIFO_WIDTH-KERNEL_SIZE;


        for (int i = 0; i <  num_additional_cycles_shifts; i++) begin
          vif.i_new_pkt <= 0;
          @(negedge vif.i_clk);
        end

      end
    end
    vif.i_new_pkt <= 0;


    for (int i = 0 ; i < 10 ; i++) begin
      $display("%d", vif.o_pixel);
      @(negedge vif.i_clk);
    end


    //`ASSERT_EQ(vif.addr, 3'b000, %3b);
    //`ASSERT_EQ(vif.payload_done, 1'b0, %b);
    @(negedge vif.i_clk);

  endtask // run

endclass // tb_cluster_kernel_size_subject_no_pad