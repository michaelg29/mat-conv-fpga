
`ifndef MAT_CONV_SVH
`define MAT_CONV_SVH

`define ACLK_PER_PS 15625 // 64MHz
`define MACCLK_PER_PS 4000  // 250MHz

`endif
