
package tb_cluster_pkg;

  import uvm_pkg::*;

  // UVM include
  `include "uvm_macros.svh"

  // utility classes
  `include "../tb_common/mat_conv.svh"
  `include "../tb_common/mat_conv_tc.svh"

  // testcases
  `include "tb_cluster_load_kernel.svh"
  `include "tb_cluster_load_kernel_block.svh"
  `include "tb_cluster_kernel_size_subject_no_pad.svh"

endpackage // tb_cluster_pkg