
package tb_input_fsm_pkg;

  import uvm_pkg::*;

  // UVM include
  `include "uvm_macros.svh"

  // utility classes
  `include "../tb_common/mat_conv.svh"
  `include "../tb_common/mat_conv_tc.svh"

  // testcases
  `include "tb_input_fsm_err_cmd.svh"
  `include "tb_input_fsm_err_proc.svh"
  `include "tb_input_fsm_valid_kern.svh"
  `include "tb_input_fsm_valid_subj.svh"

endpackage // tb_input_fsm_pkg
