class tb_global_mem_lsram_wrapper;

static task run_task();

endtask

endclass