
library ieee;
use ieee.std_logic_1164.all;

package fifo_pkg is

  

end package fifo_pkg;
