
package tb_template_pkg;

  import uvm_pkg::*;

  // UVM include
  `include "uvm_macros.svh"

  // utility classes
  `include "../tb_common/mat_conv.svh"
  `include "../tb_common/mat_conv_tc.svh"

  // testcases
  `include "tb_template_tc.svh"

endpackage // tb_template_pkg
